//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// System-Verilog Alex Grinshpun May 2018
// New coding convention dudy December 2018


module	tank_move	(	
 
					input	logic	clk,
					input	logic	resetN,
					input	logic	startOfFrame,  // short pulse every start of frame 30Hz 
					input logic collision,
					input logic [3:0] inputKeyPressed,
					output	logic	[10:0]	topLeftX,// output the top left corner 
					output	logic	[10:0]	topLeftY
					
);


// a module used to generate a ball trajectory.  

parameter int INITIAL_X = 280;
parameter int INITIAL_Y = 185;
parameter int INITIAL_X_SPEED = 0;
parameter int INITIAL_Y_SPEED = 0;
parameter int MOVEMENT_X_SPEED = 20;
parameter int MOVEMENT_Y_SPEED = 20;

const int	MULTIPLIER	=	64;
// multiplier is used to work with integers in high resolution 
// we devide at the end by multiplier which must be 2^n 
const int	x_FRAME_SIZE	=	639 * MULTIPLIER;
const int	y_FRAME_SIZE	=	479 * MULTIPLIER;


int Xspeed, topLeftX_tmp; // local parameters 
int Yspeed, topLeftY_tmp;
int flag;
int lastSpeedX;
int lastSpeedY;


//  calculation x Axis speed 

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		Xspeed	<= INITIAL_X_SPEED;
	end
	else 	begin
		if(inputKeyPressed[2] ^ inputKeyPressed[3]) begin
			if(inputKeyPressed[2]) begin
				Xspeed <= -MOVEMENT_X_SPEED;
			end
			else begin
				Xspeed <= MOVEMENT_X_SPEED;
			end
		end
		else 
			Xspeed <= 0;
	end
end


//  calculation Y Axis speed using gravity

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin 
		Yspeed	<= INITIAL_Y_SPEED;
	end 
	else 	begin
		if(inputKeyPressed[0] ^ inputKeyPressed[1]) begin
			if(inputKeyPressed[0]) begin
				Yspeed <= MOVEMENT_Y_SPEED;
			end
			else begin
				Yspeed <= -MOVEMENT_Y_SPEED;
			end
		end
		else
			Yspeed <= 0;
	end
end

// position calculate 

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN)
	begin
		topLeftX_tmp	<= INITIAL_X * MULTIPLIER;
		topLeftY_tmp	<= INITIAL_Y * MULTIPLIER;
		lastSpeedY <= INITIAL_Y_SPEED;
		lastSpeedX <= INITIAL_X_SPEED;
		flag <= 0;
	end
	else begin
		if(collision == 1'b1 && flag == 0) begin
			topLeftX_tmp  <= topLeftX_tmp - lastSpeedX; 	
			topLeftY_tmp  <= topLeftY_tmp - lastSpeedY; 
			flag <= 1;
		end
		else if (startOfFrame == 1'b1) begin // perform only 30 times per second 
				topLeftX_tmp  <= topLeftX_tmp + Xspeed; 	
				topLeftY_tmp  <= topLeftY_tmp + Yspeed; 
				lastSpeedX <= Xspeed;
				lastSpeedY <= Yspeed;
				flag <= 0;
		end
	end
end



//======--------------------------------------------------------------------------------------------------------------=
//get a better (64 times) resolution using integer   
assign 	topLeftX = topLeftX_tmp / MULTIPLIER ;   // note:  it must be 2^n 
assign 	topLeftY = topLeftY_tmp / MULTIPLIER ;    


endmodule
