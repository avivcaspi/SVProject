//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// System-Verilog Alex Grinshpun May 2018
// New coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2019 


module	brick_matrix	(	
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] pixelX,// current VGA pixel 
					input 	logic	[10:0] pixelY,
					input 	logic [10:0] topLeftX,
					input 	logic [10:0] topLeftY,
					
					output 	logic	[10:0] offsetX,// offset inside bracket from top left position 
					output 	logic	[10:0] offsetY,
					output	logic	drawingRequest, // indicates pixel inside the bracket
					output	logic	[7:0]	 RGBout, //optional color output for mux 
					output 	logic [0:13][0:16] matrix
);

parameter  int OBJECT_WIDTH_X = 544;
parameter  int OBJECT_HEIGHT_Y = 448;
parameter  logic [7:0] OBJECT_COLOR = 8'h5b ; 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// bitmap  representation for a transparent pixel 

logic [0:13][0:16] bricks_matrix = 
							'{17'b00000000000000001,
						     17'b00010100000000000,
							  17'b00010101000000000,
							  17'b00010100000000000,
							  17'b00010100000000000,
							  17'b00010100000000000,
							  17'b00100010000000000,
							  17'b00100001000000000,
							  17'b00000000000000000,
							  17'b00000000000000000,
							  17'b00000000000000000,
							  17'b00000000000000000,
							  17'b00000000000000000,
							  17'b10000000000000001};
int rightX ; //coordinates of the sides  
int bottomY ;
logic insideBracket ; 
int matrixX;
int matrixY;

//======--------------------------------------------------------------------------------------------------------------=
// Calculate object right  & bottom  boundaries
assign rightX	= (topLeftX + OBJECT_WIDTH_X);
assign bottomY	= (topLeftY + OBJECT_HEIGHT_Y);
assign matrixX = (pixelX - topLeftX) / 32;
assign matrixY = (pixelY - topLeftY) / 32;
assign matrix = bricks_matrix;

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout			<=	8'b0;
		drawingRequest	<=	1'b0;
	end
	else begin 
	
//		if ( (pixelX  >= topLeftX) &&  (pixelX < rightX) 
//			&& (pixelY  >= topLeftY) &&  (pixelY < bottomY) ) // test if it is inside the rectangle 

		//this is an example of using blocking sentence inside an always_ff block, 
		//and not waiting a clock to use the result  
		insideBracket  = 	 ( (pixelX  >= topLeftX) &&  (pixelX < rightX) // ----- LEGAL BLOCKING ASSINGMENT in ALWAYS_FF CODE 
						   && (pixelY  >= topLeftY) &&  (pixelY < bottomY) )  ; 
		
		if (insideBracket ) // test if it is inside the rectangle 
		begin 
			RGBout  <= OBJECT_COLOR ;	// colors table 
			if (bricks_matrix[matrixY][matrixX]) begin
				drawingRequest <= 1'b1;
			end
			else 
				drawingRequest <= 1'b0;
			offsetX	<= (pixelX - topLeftX) % 32; //calculate relative offsets from top left corner
			offsetY	<= (pixelY - topLeftY) % 32;
		end 
		
		else begin  
			RGBout <= TRANSPARENT_ENCODING ; // so it will not be displayed 
			drawingRequest <= 1'b0 ;// transparent color 
			offsetX	<= 0; //no offset
			offsetY	<= 0; //no offset
		end 
		
	end
end 
endmodule 