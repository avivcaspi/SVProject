

module	openBitmap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
);

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 

localparam  int OBJECT_HEIGHT_Y = 25;
localparam  int OBJECT_WIDTH_X = 100;

logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
{8'h05, 8'h29, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h29, 8'h29, 8'h04, 8'h00, 8'h29, 8'h00, 8'h00, 8'h29, 8'h00, 8'h05, 8'h29, 8'h29, 8'h04, 8'h04, 8'h29, 8'h29, 8'h29, 8'h00, 8'h05, 8'h29, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h56, 8'h5F, 8'h5F, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h5F, 8'h5F, 8'h5F, 8'h56, 8'h2D, 8'h7F, 8'h29, 8'h2D, 8'h5F, 8'h29, 8'h5A, 8'h5F, 8'h5F, 8'h32, 8'h2D, 8'h5F, 8'h5F, 8'h5F, 8'h29, 8'h56, 8'h5F, 8'h5F, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h32, 8'h56, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h5B, 8'h32, 8'h32, 8'h56, 8'h05, 8'h5F, 8'h29, 8'h05, 8'h5B, 8'h04, 8'h56, 8'h5B, 8'h5B, 8'h32, 8'h29, 8'h5B, 8'h2D, 8'h5A, 8'h29, 8'h32, 8'h56, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h00, 8'h00, 8'h29, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h2D, 8'h05, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h05, 8'h56, 8'h00, 8'h5F, 8'h29, 8'h04, 8'h56, 8'h00, 8'h56, 8'h56, 8'h32, 8'h32, 8'h04, 8'h56, 8'h00, 8'h32, 8'h29, 8'h2D, 8'h2D, 8'h25, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h2D, 8'h04, 8'h5F, 8'h56, 8'h04, 8'h56, 8'h04, 8'h2D, 8'h32, 8'h2D, 8'h2D, 8'h05, 8'h56, 8'h00, 8'h29, 8'h29, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h29, 8'h04, 8'h5B, 8'h56, 8'h04, 8'h56, 8'h04, 8'h29, 8'h32, 8'h2D, 8'h29, 8'h05, 8'h56, 8'h00, 8'h04, 8'h05, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h2D, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h29, 8'h29, 8'h00, 8'h04, 8'h56, 8'h2D, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h2D, 8'h04, 8'h00, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h05, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h2D, 8'h29, 8'h2D, 8'h04, 8'h00, 8'h05, 8'h2D, 8'h29, 8'h00, 8'h29, 8'h2D, 8'h05, 8'h00, 8'h29, 8'h2D, 8'h05, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h32, 8'h05, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h56, 8'h32, 8'h04, 8'h00, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h00, 8'h00, 8'h00, 8'h29, 8'h5F, 8'h29, 8'h00, 8'h04, 8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h2D, 8'h29, 8'h00, 8'h00, 8'h2D, 8'h2D, 8'h00, 8'h00, 8'h2D, 8'h29, 8'h29, 8'h00, 8'h29, 8'h5F, 8'h29, 8'h00, 8'h29, 8'h04, 8'h05, 8'h2D, 8'h29, 8'h29, 8'h00, 8'h29, 8'h2D, 8'h04, 8'h2D, 8'h04, 8'h00, 8'h29, 8'h2D, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h2D, 8'h32, 8'h04, 8'h5F, 8'h56, 8'h5F, 8'h2D, 8'h00, 8'h32, 8'h5F, 8'h56, 8'h00, 8'h56, 8'h5B, 8'h32, 8'h04, 8'h5A, 8'h5A, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h56, 8'h29, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h5A, 8'h5A, 8'h04, 8'h00, 8'h2D, 8'h32, 8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h5F, 8'h32, 8'h00, 8'h29, 8'h5F, 8'h5B, 8'h04, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h5F, 8'h5A, 8'h00, 8'h04, 8'h5F, 8'h5F, 8'h05, 8'h04, 8'h5F, 8'h56, 8'h5B, 8'h00, 8'h2D, 8'h5F, 8'h52, 8'h00, 8'h32, 8'h29, 8'h2D, 8'h5B, 8'h56, 8'h56, 8'h00, 8'h56, 8'h5F, 8'h05, 8'h5F, 8'h29, 8'h00, 8'h56, 8'h5F, 8'h32, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h5B, 8'h5B, 8'h29, 8'h00, 8'h56, 8'h5B, 8'h32, 8'h32, 8'h00, 8'h56, 8'h2D, 8'h56, 8'h05, 8'h56, 8'h2D, 8'h56, 8'h05, 8'h56, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h5F, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h2D, 8'h29, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h5F, 8'h5B, 8'h04, 8'h00, 8'h2D, 8'h5B, 8'h5B, 8'h29, 8'h00, 8'h00, 8'h00, 8'h29, 8'h5B, 8'h05, 8'h00, 8'h32, 8'h2D, 8'h32, 8'h29, 8'h00, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h56, 8'h04, 8'h29, 8'h32, 8'h32, 8'h2D, 8'h00, 8'h5A, 8'h32, 8'h56, 8'h05, 8'h04, 8'h5B, 8'h05, 8'h00, 8'h32, 8'h29, 8'h04, 8'h5B, 8'h2D, 8'h56, 8'h00, 8'h2D, 8'h56, 8'h00, 8'h56, 8'h29, 8'h00, 8'h56, 8'h2D, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h5B, 8'h56, 8'h04, 8'h00, 8'h56, 8'h5B, 8'h29, 8'h56, 8'h05, 8'h56, 8'h00, 8'h56, 8'h29, 8'h56, 8'h04, 8'h32, 8'h29, 8'h56, 8'h04, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h5F, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h29, 8'h2D, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h5F, 8'h5B, 8'h04, 8'h00, 8'h2D, 8'h5B, 8'h5A, 8'h29, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h56, 8'h04, 8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h00, 8'h2D, 8'h05, 8'h32, 8'h29, 8'h05, 8'h56, 8'h00, 8'h56, 8'h2D, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h5B, 8'h29, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h29, 8'h29, 8'h32, 8'h00, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h2D, 8'h5A, 8'h2D, 8'h32, 8'h00, 8'h56, 8'h29, 8'h5F, 8'h05, 8'h29, 8'h29, 8'h5F, 8'h00, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h2D, 8'h56, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h56, 8'h04, 8'h00, 8'h2D, 8'h32, 8'h29, 8'h32, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h05, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h00, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h04, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h2D, 8'h00, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h29, 8'h2D, 8'h2D, 8'h56, 8'h32, 8'h56, 8'h04, 8'h56, 8'h56, 8'h2D, 8'h04, 8'h5B, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h05, 8'h32, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h32, 8'h04, 8'h00, 8'h2D, 8'h2D, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h04, 8'h56, 8'h04, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h56, 8'h32, 8'h32, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h2D, 8'h5F, 8'h5F, 8'h32, 8'h00, 8'h32, 8'h83, 8'h32, 8'h00, 8'h56, 8'h83, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h29, 8'h29, 8'h00, 8'h04, 8'h56, 8'h00, 8'h32, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h56, 8'h29, 8'h04, 8'h00, 8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h04, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h5F, 8'h5F, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h2D, 8'h56, 8'h29, 8'h04, 8'h04, 8'h2D, 8'h32, 8'h5A, 8'h04, 8'h29, 8'h56, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h29, 8'h04, 8'h56, 8'h00, 8'h56, 8'h5A, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h56, 8'h04, 8'h04, 8'h04, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h04, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h32, 8'h29, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h29, 8'h32, 8'h00, 8'h04, 8'h05, 8'h2D, 8'h05, 8'h5B, 8'h29, 8'h29, 8'h29, 8'h5B, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h2D, 8'h04, 8'h56, 8'h00, 8'h56, 8'h5B, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h00, 8'h29, 8'h29, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h04, 8'h04, 8'h56, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h00, 8'h56, 8'h05, 8'h04, 8'h56, 8'h00, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h04, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h56, 8'h00, 8'h56, 8'h05, 8'h2D, 8'h2D, 8'h00, 8'h04, 8'h00, 8'h04, 8'h04, 8'h04, 8'h05, 8'h00 },
{8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h32, 8'h29, 8'h56, 8'h00, 8'h56, 8'h29, 8'h32, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h04, 8'h52, 8'h04, 8'h56, 8'h00, 8'h32, 8'h5B, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h00, 8'h2D, 8'h29, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h05, 8'h56, 8'h29, 8'h04, 8'h56, 8'h04, 8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h00, 8'h2D, 8'h29, 8'h32, 8'h29, 8'h29, 8'h32, 8'h00, 8'h56, 8'h04, 8'h32, 8'h29, 8'h04, 8'h56, 8'h29, 8'h04, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h00, 8'h29, 8'h5B, 8'h04, 8'h5F, 8'h05, 8'h05, 8'h56, 8'h00, 8'h32, 8'h29, 8'h2D, 8'h2D, 8'h29, 8'h32, 8'h04 },
{8'h32, 8'h56, 8'h00, 8'h00, 8'h00, 8'h5B, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h32, 8'h56, 8'h56, 8'h05, 8'h56, 8'h32, 8'h32, 8'h29, 8'h32, 8'h32, 8'h32, 8'h00, 8'h00, 8'h04, 8'h5B, 8'h56, 8'h56, 8'h56, 8'h29, 8'h5B, 8'h04, 8'h2D, 8'h5F, 8'h04, 8'h00, 8'h56, 8'h32, 8'h00, 8'h2D, 8'h5B, 8'h32, 8'h5B, 8'h29, 8'h32, 8'h56, 8'h04, 8'h5B, 8'h29, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h00, 8'h2D, 8'h56, 8'h56, 8'h05, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h56, 8'h56, 8'h04, 8'h29, 8'h56, 8'h56, 8'h29, 8'h00, 8'h5B, 8'h29, 8'h32, 8'h32, 8'h00, 8'h56, 8'h32, 8'h04, 8'h56, 8'h32, 8'h29, 8'h5F, 8'h29, 8'h56, 8'h29, 8'h04, 8'h5B, 8'h56, 8'h5B, 8'h2D, 8'h00, 8'h56, 8'h56, 8'h32, 8'h29, 8'h32, 8'h2E, 8'h2D, 8'h56, 8'h04 },
{8'h5B, 8'h5F, 8'h00, 8'h00, 8'h04, 8'h7F, 8'h56, 8'h00, 8'h00, 8'h00, 8'h32, 8'h83, 8'h56, 8'h04, 8'h32, 8'h7F, 8'h32, 8'h04, 8'h32, 8'h83, 8'h2D, 8'h00, 8'h00, 8'h05, 8'h7F, 8'h5F, 8'h83, 8'h56, 8'h2D, 8'h83, 8'h29, 8'h2D, 8'h83, 8'h29, 8'h00, 8'h5F, 8'h56, 8'h00, 8'h32, 8'h83, 8'h5F, 8'h83, 8'h29, 8'h5A, 8'h5B, 8'h29, 8'h83, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h00, 8'h29, 8'h83, 8'h5F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h83, 8'h5B, 8'h00, 8'h04, 8'h5F, 8'h5F, 8'h04, 8'h05, 8'h83, 8'h32, 8'h32, 8'h5A, 8'h00, 8'h52, 8'h56, 8'h00, 8'h5F, 8'h56, 8'h2D, 8'h83, 8'h29, 8'h5B, 8'h32, 8'h00, 8'h5B, 8'h5B, 8'h5A, 8'h56, 8'h00, 8'h56, 8'h83, 8'h32, 8'h29, 8'h32, 8'h32, 8'h2D, 8'h56, 8'h04 },
{8'h04, 8'h05, 8'h00, 8'h00, 8'h00, 8'h05, 8'h04, 8'h00, 8'h00, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h00, 8'h00, 8'h05, 8'h05, 8'h05, 8'h04, 8'h04, 8'h05, 8'h00, 8'h04, 8'h05, 8'h00, 8'h00, 8'h05, 8'h04, 8'h00, 8'h04, 8'h05, 8'h05, 8'h05, 8'h00, 8'h04, 8'h04, 8'h00, 8'h05, 8'h04, 8'h00, 8'h00, 8'h00, 8'h04, 8'h04, 8'h00, 8'h00, 8'h05, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h04, 8'h00, 8'h00, 8'h05, 8'h05, 8'h00, 8'h00, 8'h05, 8'h04, 8'h04, 8'h04, 8'h00, 8'h04, 8'h04, 8'h00, 8'h05, 8'h04, 8'h04, 8'h05, 8'h00, 8'h04, 8'h04, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 }
};

// pipeline (ff) to get the pixel color from the array 	 

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1 )  // inside an external bracket 
			RGBout <= object_colors[offsetY][offsetX];	//get RGB from the colors table  
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end

//======--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule