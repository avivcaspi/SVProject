const logic [0:13] [0:16] [2:0] map1 = {
{3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h4, 3'h3, 3'h3, 3'h3, 3'h4, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h4, 3'h4, 3'h4, 3'h4, 3'h4, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h4, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h3, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h0, 3'h0, 3'h4 },
{3'h0, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h3, 3'h3, 3'h0, 3'h0 },
{3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h3, 3'h3, 3'h4, 3'h0, 3'h3, 3'h4, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h4, 3'h3, 3'h3, 3'h4, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0 }};

const logic [0:13] [0:16] [2:0] map2 = {
{3'h0, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h4, 3'h4, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h3, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h4, 3'h0, 3'h4, 3'h3, 3'h0, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0 },
{3'h4, 3'h0, 3'h0, 3'h3, 3'h0, 3'h4, 3'h4, 3'h3, 3'h4, 3'h4, 3'h3, 3'h4, 3'h0, 3'h3, 3'h0, 3'h0, 3'h4 },
{3'h4, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h4 },
{3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h0, 3'h4, 3'h4, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h3, 3'h3, 3'h4, 3'h4, 3'h0, 3'h0, 3'h0 },
{3'h4, 3'h3, 3'h0, 3'h4, 3'h4, 3'h3, 3'h3, 3'h3, 3'h0, 3'h0, 3'h3, 3'h3, 3'h4, 3'h4, 3'h0, 3'h3, 3'h4 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h4, 3'h4, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h4, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h3, 3'h4, 3'h0, 3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0 }};


const logic [0:13] [0:16] [2:0] map3 = {
{3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0 },
{3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h3, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h3, 3'h4, 3'h4, 3'h4, 3'h0, 3'h4, 3'h4, 3'h4, 3'h4, 3'h0, 3'h4, 3'h4, 3'h4, 3'h4, 3'h4 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h3, 3'h0, 3'h4, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h4, 3'h0, 3'h3, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h3, 3'h4, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h4, 3'h0, 3'h3, 3'h3, 3'h0, 3'h0, 3'h3, 3'h3, 3'h3, 3'h0, 3'h4, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h3, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h0, 3'h4, 3'h0, 3'h3, 3'h4, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0, 3'h3, 3'h4, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h3, 3'h0, 3'h4, 3'h0, 3'h0, 3'h4, 3'h3, 3'h0, 3'h4, 3'h3, 3'h0, 3'h3, 3'h4, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h3, 3'h4, 3'h4, 3'h4, 3'h0, 3'h4, 3'h4, 3'h4, 3'h4, 3'h0, 3'h0, 3'h0, 3'h4, 3'h0, 3'h0 },
{3'h0, 3'h3, 3'h3, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h4, 3'h3, 3'h0 },
{3'h0, 3'h3, 3'h0, 3'h3, 3'h0, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h3, 3'h0, 3'h3, 3'h0 },
{3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0, 3'h0}};