localparam  int OBJECT_HEIGHT_Y = 32;
localparam  int OBJECT_WIDTH_X = 32;

logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'hB6, 8'hDB, 8'h6D, 8'h24, 8'h24, 8'h6D, 8'hDB, 8'hB6, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hDB, 8'hB6, 8'h24, 8'h49, 8'hDB, 8'hDB, 8'h49, 8'h24, 8'hB6, 8'hDB, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'hDA, 8'hDB, 8'h49, 8'h24, 8'hB6, 8'hFF, 8'h92, 8'h92, 8'hFF, 8'hB6, 8'h24, 8'h49, 8'hDB, 8'hDA, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h92, 8'hFF, 8'h92, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'h49, 8'h25, 8'h25, 8'h49, 8'hFF, 8'hFF, 8'h6D, 8'h00, 8'h92, 8'hFF, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hDB, 8'hB6, 8'h24, 8'h25, 8'hDA, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'hFF, 8'hFF, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hDA, 8'h25, 8'h24, 8'hB6, 8'hDB, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h24, 8'hB6, 8'hDB, 8'h6D, 8'h24, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h24, 8'h92, 8'h92, 8'h24, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h24, 8'h6D, 8'hDB, 8'hB6, 8'h24, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h92, 8'hFF, 8'h92, 8'h24, 8'h49, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h49, 8'h49, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h49, 8'h24, 8'h92, 8'hFF, 8'h92, 8'h00, 8'h00 },
{8'h00, 8'h49, 8'hDA, 8'h49, 8'h24, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h24, 8'h49, 8'hDA, 8'h49, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h92, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'h92, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h25, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h25, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h24, 8'h92, 8'h92, 8'h92, 8'h92, 8'h00, 8'h92, 8'h92, 8'h92, 8'hB6, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'hB6, 8'h92, 8'h92, 8'h92, 8'h00, 8'h92, 8'h92, 8'h92, 8'h92, 8'h24, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h24, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h00, 8'h6D, 8'h6D, 8'h6D, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'h123, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'h123, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'h123, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'h123, 8'hDB, 8'h00, 8'h00, 8'h00, 8'hDB, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h92, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h92, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h6D, 8'h92, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h24, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h00, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h6D, 8'h6D, 8'h6D, 8'h49, 8'h00, 8'h49, 8'h6D, 8'h6D, 8'h6D, 8'h24, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h24, 8'hB6, 8'hB6, 8'hB6, 8'h92, 8'h00, 8'h92, 8'hB6, 8'hB6, 8'hB6, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'hB6, 8'hB6, 8'hB6, 8'h92, 8'h00, 8'h92, 8'hB6, 8'hB6, 8'hB6, 8'h24, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h49, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'h49, 8'h00, 8'h00 },
{8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00 },
{8'h00, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hB6, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 }
};

wire [7:0] red_sig, green_sig, blue_sig;
assign red_sig     = {object_colors[offsetY][offsetX][7:5] , 5'd0};
assign green_sig   = {object_colors[offsetY][offsetX][4:2] , 5'd0};
assign blue_sig    = {object_colors[offsetY][offsetX][1:0] , 6'd0};


