localparam  int OBJECT_HEIGHT_Y = 25;
localparam  int OBJECT_WIDTH_X = 100;

logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {
{8'h05, 8'h29, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h29, 8'h29, 8'h04, 8'h00, 8'h29, 8'h00, 8'h00, 8'h29, 8'h00, 8'h05, 8'h29, 8'h29, 8'h04, 8'h04, 8'h29, 8'h29, 8'h29, 8'h00, 8'h05, 8'h29, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h56, 8'h5F, 8'h5F, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h5F, 8'h5F, 8'h5F, 8'h56, 8'h2D, 8'h7F, 8'h29, 8'h2D, 8'h5F, 8'h29, 8'h5A, 8'h5F, 8'h5F, 8'h32, 8'h2D, 8'h5F, 8'h5F, 8'h5F, 8'h29, 8'h56, 8'h5F, 8'h5F, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h32, 8'h56, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h5B, 8'h32, 8'h32, 8'h56, 8'h05, 8'h5F, 8'h29, 8'h05, 8'h5B, 8'h04, 8'h56, 8'h5B, 8'h5B, 8'h32, 8'h29, 8'h5B, 8'h2D, 8'h5A, 8'h29, 8'h32, 8'h56, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h00, 8'h00, 8'h29, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h2D, 8'h05, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h05, 8'h56, 8'h00, 8'h5F, 8'h29, 8'h04, 8'h56, 8'h00, 8'h56, 8'h56, 8'h32, 8'h32, 8'h04, 8'h56, 8'h00, 8'h32, 8'h29, 8'h2D, 8'h2D, 8'h25, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h2D, 8'h04, 8'h5F, 8'h56, 8'h04, 8'h56, 8'h04, 8'h2D, 8'h32, 8'h2D, 8'h2D, 8'h05, 8'h56, 8'h00, 8'h29, 8'h29, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h29, 8'h04, 8'h5B, 8'h56, 8'h04, 8'h56, 8'h04, 8'h29, 8'h32, 8'h2D, 8'h29, 8'h05, 8'h56, 8'h00, 8'h04, 8'h05, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h2D, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h29, 8'h29, 8'h00, 8'h04, 8'h56, 8'h2D, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h2D, 8'h04, 8'h00, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h05, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h2D, 8'h29, 8'h2D, 8'h04, 8'h00, 8'h05, 8'h2D, 8'h29, 8'h00, 8'h29, 8'h2D, 8'h05, 8'h00, 8'h29, 8'h2D, 8'h05, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h32, 8'h05, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h56, 8'h32, 8'h04, 8'h00, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h00, 8'h00, 8'h00, 8'h29, 8'h5F, 8'h29, 8'h00, 8'h04, 8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h2D, 8'h29, 8'h00, 8'h00, 8'h2D, 8'h2D, 8'h00, 8'h00, 8'h2D, 8'h29, 8'h29, 8'h00, 8'h29, 8'h5F, 8'h29, 8'h00, 8'h29, 8'h04, 8'h05, 8'h2D, 8'h29, 8'h29, 8'h00, 8'h29, 8'h2D, 8'h04, 8'h2D, 8'h04, 8'h00, 8'h29, 8'h2D, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h2D, 8'h32, 8'h04, 8'h5F, 8'h56, 8'h5F, 8'h2D, 8'h00, 8'h32, 8'h5F, 8'h56, 8'h00, 8'h56, 8'h5B, 8'h32, 8'h04, 8'h5A, 8'h5A, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h56, 8'h29, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h5A, 8'h5A, 8'h04, 8'h00, 8'h2D, 8'h32, 8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h5F, 8'h32, 8'h00, 8'h29, 8'h5F, 8'h5B, 8'h04, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h5F, 8'h5A, 8'h00, 8'h04, 8'h5F, 8'h5F, 8'h05, 8'h04, 8'h5F, 8'h56, 8'h5B, 8'h00, 8'h2D, 8'h5F, 8'h52, 8'h00, 8'h32, 8'h29, 8'h2D, 8'h5B, 8'h56, 8'h56, 8'h00, 8'h56, 8'h5F, 8'h05, 8'h5F, 8'h29, 8'h00, 8'h56, 8'h5F, 8'h32, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h5B, 8'h5B, 8'h29, 8'h00, 8'h56, 8'h5B, 8'h32, 8'h32, 8'h00, 8'h56, 8'h2D, 8'h56, 8'h05, 8'h56, 8'h2D, 8'h56, 8'h05, 8'h56, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h5F, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h2D, 8'h29, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h5F, 8'h5B, 8'h04, 8'h00, 8'h2D, 8'h5B, 8'h5B, 8'h29, 8'h00, 8'h00, 8'h00, 8'h29, 8'h5B, 8'h05, 8'h00, 8'h32, 8'h2D, 8'h32, 8'h29, 8'h00, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h56, 8'h04, 8'h29, 8'h32, 8'h32, 8'h2D, 8'h00, 8'h5A, 8'h32, 8'h56, 8'h05, 8'h04, 8'h5B, 8'h05, 8'h00, 8'h32, 8'h29, 8'h04, 8'h5B, 8'h2D, 8'h56, 8'h00, 8'h2D, 8'h56, 8'h00, 8'h56, 8'h29, 8'h00, 8'h56, 8'h2D, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h5B, 8'h56, 8'h04, 8'h00, 8'h56, 8'h5B, 8'h29, 8'h56, 8'h05, 8'h56, 8'h00, 8'h56, 8'h29, 8'h56, 8'h04, 8'h32, 8'h29, 8'h56, 8'h04, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h5F, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h29, 8'h2D, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h5F, 8'h5B, 8'h04, 8'h00, 8'h2D, 8'h5B, 8'h5A, 8'h29, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h56, 8'h04, 8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h00, 8'h2D, 8'h05, 8'h32, 8'h29, 8'h05, 8'h56, 8'h00, 8'h56, 8'h2D, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h5B, 8'h29, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h29, 8'h29, 8'h32, 8'h00, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h2D, 8'h5A, 8'h2D, 8'h32, 8'h00, 8'h56, 8'h29, 8'h5F, 8'h05, 8'h29, 8'h29, 8'h5F, 8'h00, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h2D, 8'h56, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h56, 8'h04, 8'h00, 8'h2D, 8'h32, 8'h29, 8'h32, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h05, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h00, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h04, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h2D, 8'h00, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h29, 8'h2D, 8'h2D, 8'h56, 8'h32, 8'h56, 8'h04, 8'h56, 8'h56, 8'h2D, 8'h04, 8'h5B, 8'h32, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h2D, 8'h00, 8'h04, 8'h56, 8'h05, 8'h32, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h32, 8'h04, 8'h00, 8'h2D, 8'h2D, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h04, 8'h56, 8'h04, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h56, 8'h32, 8'h32, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h2D, 8'h5F, 8'h5F, 8'h32, 8'h00, 8'h32, 8'h83, 8'h32, 8'h00, 8'h56, 8'h83, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h29, 8'h29, 8'h00, 8'h04, 8'h56, 8'h00, 8'h32, 8'h56, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h56, 8'h29, 8'h04, 8'h00, 8'h2D, 8'h32, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h04, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h5F, 8'h5F, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h2D, 8'h56, 8'h29, 8'h04, 8'h04, 8'h2D, 8'h32, 8'h5A, 8'h04, 8'h29, 8'h56, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h29, 8'h04, 8'h56, 8'h00, 8'h56, 8'h5A, 8'h00, 8'h00, 8'h32, 8'h2D, 8'h00, 8'h05, 8'h56, 8'h04, 8'h04, 8'h04, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h56, 8'h00, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h00, 8'h56, 8'h04, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h32, 8'h00, 8'h56, 8'h05, 8'h32, 8'h32, 8'h29, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h2D, 8'h32, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h29, 8'h32, 8'h00, 8'h04, 8'h05, 8'h2D, 8'h05, 8'h5B, 8'h29, 8'h29, 8'h29, 8'h5B, 8'h00, 8'h00, 8'h00, 8'h56, 8'h05, 8'h00, 8'h2D, 8'h04, 8'h56, 8'h00, 8'h56, 8'h5B, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h00, 8'h29, 8'h29, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h04, 8'h56, 8'h04, 8'h04, 8'h56, 8'h00, 8'h29, 8'h56, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h04, 8'h00, 8'h56, 8'h05, 8'h04, 8'h56, 8'h00, 8'h56, 8'h05, 8'h32, 8'h29, 8'h04, 8'h56, 8'h04, 8'h00, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h04, 8'h29, 8'h56, 8'h00, 8'h56, 8'h05, 8'h2D, 8'h2D, 8'h00, 8'h04, 8'h00, 8'h04, 8'h04, 8'h04, 8'h05, 8'h00 },
{8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h00, 8'h04, 8'h56, 8'h00, 8'h32, 8'h29, 8'h56, 8'h00, 8'h56, 8'h29, 8'h32, 8'h04, 8'h56, 8'h00, 8'h00, 8'h00, 8'h56, 8'h04, 8'h04, 8'h52, 8'h04, 8'h56, 8'h00, 8'h32, 8'h5B, 8'h00, 8'h00, 8'h32, 8'h29, 8'h00, 8'h05, 8'h56, 8'h00, 8'h2D, 8'h29, 8'h2D, 8'h2D, 8'h00, 8'h56, 8'h04, 8'h00, 8'h00, 8'h05, 8'h56, 8'h29, 8'h04, 8'h56, 8'h04, 8'h2D, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h00, 8'h2D, 8'h29, 8'h32, 8'h29, 8'h29, 8'h32, 8'h00, 8'h56, 8'h04, 8'h32, 8'h29, 8'h04, 8'h56, 8'h29, 8'h04, 8'h32, 8'h29, 8'h00, 8'h56, 8'h00, 8'h56, 8'h00, 8'h29, 8'h5B, 8'h04, 8'h5F, 8'h05, 8'h05, 8'h56, 8'h00, 8'h32, 8'h29, 8'h2D, 8'h2D, 8'h29, 8'h32, 8'h04 },
{8'h32, 8'h56, 8'h00, 8'h00, 8'h00, 8'h5B, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h32, 8'h56, 8'h56, 8'h05, 8'h56, 8'h32, 8'h32, 8'h29, 8'h32, 8'h32, 8'h32, 8'h00, 8'h00, 8'h04, 8'h5B, 8'h56, 8'h56, 8'h56, 8'h29, 8'h5B, 8'h04, 8'h2D, 8'h5F, 8'h04, 8'h00, 8'h56, 8'h32, 8'h00, 8'h2D, 8'h5B, 8'h32, 8'h5B, 8'h29, 8'h32, 8'h56, 8'h04, 8'h5B, 8'h29, 8'h00, 8'h00, 8'h00, 8'h56, 8'h2D, 8'h00, 8'h2D, 8'h56, 8'h56, 8'h05, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h56, 8'h56, 8'h04, 8'h29, 8'h56, 8'h56, 8'h29, 8'h00, 8'h5B, 8'h29, 8'h32, 8'h32, 8'h00, 8'h56, 8'h32, 8'h04, 8'h56, 8'h32, 8'h29, 8'h5F, 8'h29, 8'h56, 8'h29, 8'h04, 8'h5B, 8'h56, 8'h5B, 8'h2D, 8'h00, 8'h56, 8'h56, 8'h32, 8'h29, 8'h32, 8'h2E, 8'h2D, 8'h56, 8'h04 },
{8'h5B, 8'h5F, 8'h00, 8'h00, 8'h04, 8'h7F, 8'h56, 8'h00, 8'h00, 8'h00, 8'h32, 8'h83, 8'h56, 8'h04, 8'h32, 8'h7F, 8'h32, 8'h04, 8'h32, 8'h83, 8'h2D, 8'h00, 8'h00, 8'h05, 8'h7F, 8'h5F, 8'h83, 8'h56, 8'h2D, 8'h83, 8'h29, 8'h2D, 8'h83, 8'h29, 8'h00, 8'h5F, 8'h56, 8'h00, 8'h32, 8'h83, 8'h5F, 8'h83, 8'h29, 8'h5A, 8'h5B, 8'h29, 8'h83, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h56, 8'h56, 8'h00, 8'h29, 8'h83, 8'h5F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h83, 8'h5B, 8'h00, 8'h04, 8'h5F, 8'h5F, 8'h04, 8'h05, 8'h83, 8'h32, 8'h32, 8'h5A, 8'h00, 8'h52, 8'h56, 8'h00, 8'h5F, 8'h56, 8'h2D, 8'h83, 8'h29, 8'h5B, 8'h32, 8'h00, 8'h5B, 8'h5B, 8'h5A, 8'h56, 8'h00, 8'h56, 8'h83, 8'h32, 8'h29, 8'h32, 8'h32, 8'h2D, 8'h56, 8'h04 },
{8'h04, 8'h05, 8'h00, 8'h00, 8'h00, 8'h05, 8'h04, 8'h00, 8'h00, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h00, 8'h00, 8'h05, 8'h05, 8'h05, 8'h04, 8'h04, 8'h05, 8'h00, 8'h04, 8'h05, 8'h00, 8'h00, 8'h05, 8'h04, 8'h00, 8'h04, 8'h05, 8'h05, 8'h05, 8'h00, 8'h04, 8'h04, 8'h00, 8'h05, 8'h04, 8'h00, 8'h00, 8'h00, 8'h04, 8'h04, 8'h00, 8'h00, 8'h05, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h04, 8'h00, 8'h00, 8'h05, 8'h05, 8'h00, 8'h00, 8'h05, 8'h04, 8'h04, 8'h04, 8'h00, 8'h04, 8'h04, 8'h00, 8'h05, 8'h04, 8'h04, 8'h05, 8'h00, 8'h04, 8'h04, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00, 8'h04, 8'h05, 8'h04, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 },
{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00 }
};

wire [7:0] red_sig, green_sig, blue_sig;
assign red_sig     = {object_colors[offsetY][offsetX][7:5] , 5'd0};
assign green_sig   = {object_colors[offsetY][offsetX][4:2] , 5'd0};
assign blue_sig    = {object_colors[offsetY][offsetX][1:0] , 6'd0};


